class adder_trans;
  
  randc logic [3:0]  a_i;
  randc logic [3:0]  b_i;
        logic [4:0]  s_o;

endclass