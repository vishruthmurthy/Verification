module environment();

and_2_if and_2_intf ();

driver drv (and_2_intf);
monitor mon (and_2_intf);
scoreboard sb (and_2_intf);

endmodule
