class counter_trans;
  
  randc logic       enable_i;
  randc logic       load_i;
  randc logic [3:0] data_i;
        logic [3:0] count_o;

endclass