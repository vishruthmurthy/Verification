module adder (
	input [3:0] a,
	input [3:0] b,
	output [4:0] s
	);

assign s= a+b;

endmodule
