//---------------------------------------------------------------------------
// Title       : 4-Bit Adder Simple Verification Environment
// Design      : Driver
// File        : driver.sv
//---------------------------------------------------------------------------

class driver;

  virtual adder_if.drv_mp drv_if;
  
  // Override the constructor to connect with interface
  function new(virtual adder_if.drv_mp intf);
    drv_if = intf;
  endfunction
  
  // Task to drive input signals of interface
  // Get the values for A and B generated by generator
  task drive(input logic [3:0] a, input logic [3:0] b);
    drv_if.a = a;
    drv_if.b = b;
    $display($time, "ns [DRV] : A = %d, B = %d", drv_if.a, drv_if.b);
  endtask
  
endclass